`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:33:54 04/26/2017 
// Design Name: 
// Module Name:    cordic 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module cordic(
    input [32:0] x_in,
    input [32:0] k_in,
    input [32:0] y_in,
    input [32:0] e_k_in,
    input CE,
    output [32:0] n_out,
    output done,
    output [32:0] y_out
    );


endmodule
